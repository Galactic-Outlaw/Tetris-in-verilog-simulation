
module tetris1_testmodule();
reg Reset,Clk,Start,try_again,Left,Right,Down,Rotate;
wire [159:0] blocks;
wire [7:0] score;
wire [1:0] orientation;
wire [7:0] position;
wire [2:0] next_block;
wire O_Initial,O_Generate,O_Rotate,O_Collision,O_Lose;

tetris1 test( Reset, Clk, Start, try_again, Left, Right, Down, Rotate,
	O_Initial, O_Generate, O_Rotate, O_Collision, O_Lose, blocks, score, orientation, position, next_block
    );
initial
begin
$dumpfile("demo_test.vcd");
$dumpvars(0,tetris1_testmodule);
end
initial
begin
Reset=1;
Clk=0;
Start=0;
try_again=0;
Left=0;
Right=0;
Down=0;
Rotate=0;
#10;
Reset=0;
Clk=1;
Start=1;
try_again=0;
Left=0;
Right=0;
Down=0;
Rotate=0;
#10;
Reset=0;
Clk=0;
Start=0;
try_again=0;
Left=0;
Right=0;
Down=0;
Rotate=0;
#10;
Reset=0;
Clk=1;
Start=0;
try_again=0;
Left=0;
Right=0;
Down=0;
Rotate=1;
#10;
Reset=0;
Clk=0;
Start=0;
try_again=0;
Left=0;
Right=0;
Down=0;
Rotate=0;
#10;
Reset=0;
Clk=1;
Start=0;
try_again=0;
Left=0;
Right=0;
Down=1;
Rotate=0;
#10;
Reset=0;
Clk=0;
Start=0;
try_again=0;
Left=0;
Right=0;
Down=0;
Rotate=0;
#10;
Reset=0;
Clk=1;
Start=0;
try_again=0;
Left=0;
Right=0;
Down=1;
Rotate=0;
#10;
Reset=0;
Clk=0;
Start=0;
try_again=0;
Left=0;
Right=0;
Down=0;
Rotate=0;
#10;
Reset=0;
Clk=1;
Start=0;
try_again=0;
Left=0;
Right=0;
Down=1;
Rotate=0;
#10;
Reset=0;
Clk=0;
Start=0;
try_again=0;
Left=0;
Right=0;
Down=0;
Rotate=0;
#10;
Reset=0;
Clk=1;
Start=0;
try_again=0;
Left=0;
Right=1;
Down=0;
Rotate=0;
#10;
Reset=0;
Clk=0;
Start=0;
try_again=0;
Left=0;
Right=0;
Down=0;
Rotate=0;
#10;
Reset=0;
Clk=1;
Start=0;
try_again=0;
Left=1;
Right=0;
Down=0;
Rotate=0;
#10;
end
endmodule
